module Adder(
    input wire [31:0] operandA, // 피연산자 A
    input wire [31:0] operandB, // 피연산자 B
    output reg [31:0] sum       // 덧셈 결과
);

    always @* begin
        // 두 피연산자를 더하기
        sum = operandA + operandB;
    end

endmodule
