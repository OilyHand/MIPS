module WB_Stage(
    input [31:0] MEMtoWB_ReadData,
    input [31:0] MEMtoWB_ALU_result,
// need to add control signals
    output [31:0] WB_WriteData,
    output [31:0] WB_RegDest
    );
    // MUX
    
endmodule
