module MEM_Stage(
    input [31:0] EXtoMEM_ALU_result,
    input [31:0] EXtoMEM_RegDest,
// need to add control signals
    output [31:0] ReadData,
    output [31:0] MEMtoWB_ALU_result,
    output [31:0] MEMtoWB_RegDest
    );
    // Data Memory
endmodule
